module filelock

// TODO : implement

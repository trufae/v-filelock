module filelock

// TODO

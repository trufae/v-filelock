module filelock

// TODO: move the current code in lib.v into here
